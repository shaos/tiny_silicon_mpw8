module gpio_defaults_block_0c00 (VGND,
    VPWR,
    gpio_defaults);
 input VGND;
 input VPWR;
 output [12:0] gpio_defaults;

 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;
 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[1] ;

 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign gpio_defaults[0] = \gpio_defaults_low[0] ;
 assign gpio_defaults[1] = \gpio_defaults_low[1] ;
 assign gpio_defaults[2] = \gpio_defaults_low[2] ;
 assign gpio_defaults[3] = \gpio_defaults_low[3] ;
 assign gpio_defaults[4] = \gpio_defaults_low[4] ;
 assign gpio_defaults[5] = \gpio_defaults_low[5] ;
 assign gpio_defaults[6] = \gpio_defaults_low[6] ;
 assign gpio_defaults[7] = \gpio_defaults_low[7] ;
 assign gpio_defaults[8] = \gpio_defaults_low[8] ;
 assign gpio_defaults[9] = \gpio_defaults_low[9] ;
 assign gpio_defaults[10] = \gpio_defaults_high[10] ;
 assign gpio_defaults[11] = \gpio_defaults_high[11] ;
 assign gpio_defaults[12] = \gpio_defaults_low[12] ;
endmodule
